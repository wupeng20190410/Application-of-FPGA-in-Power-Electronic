module (
        input           wire            a,
        input           wire            b

)


endmodule