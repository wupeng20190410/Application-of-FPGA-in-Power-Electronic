module (
        input           wire           d,
        input           wire            fg,
        output          reg             c

)

assign c = a |b;


endmodule