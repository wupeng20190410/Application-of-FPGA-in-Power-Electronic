module (
        input           wire            a,
        input           wire            b,
        output          reg             c

)

always @() begin
        
end


endmodule