module adder (
        input           wire            a,
        input           wire            b,
        output          reg             c

)
assign c = a & b;



endmodule